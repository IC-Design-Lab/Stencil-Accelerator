reg [`BW-1:0] golden_item0   ;    
reg [`BW-1:0] golden_item1   ;    
reg [`BW-1:0] golden_item2   ;    
reg [`BW-1:0] dut_item0      ;    
reg [`BW-1:0] dut_item1      ;    
reg [`BW-1:0] dut_item2      ;    

real golden_real_item0   ;  
real golden_real_item1   ;  
real golden_real_item2   ;  
real dut_real_item0      ;
real dut_real_item1      ;
real dut_real_item2      ;

real error_percent0   ;    
real error_percent1   ;    
real error_percent2   ;    

